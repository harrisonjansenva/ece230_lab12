// Implement binary state machine
module binary (
    input w,
    input clk,
    input reset,
    output z,
    output [3:0] state
);
wire Anext, Bnext, Cnext, Dnext;


endmodule

